LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ALU_TB IS
-- empty
END ENTITY;

ARCHITECTURE TB_ARCH OF ALU_TB IS

SIGNAL A : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
SIGNAL B : STD_LOGIC_VECTOR(7 DOWNTO 0) := "00000000";
SIGNAL CONTROL_BUS : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
SIGNAL Y : STD_LOGIC_VECTOR(7 DOWNTO 0);

-- DUT component
COMPONENT ALU IS
  PORT(
    a: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    b: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    control_bus: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
    y: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
  );
END COMPONENT;

BEGIN

  -- Connect DUT
  UUT: ALU PORT MAP(A, B, CONTROL_BUS, Y);

  PROCESS
  BEGIN
    -- Test case 1: A AND B
    A <= X"0A";
    B <= X"0B";
    CONTROL_BUS <= "000";
    WAIT FOR 100 ns;
    
    assert false report "Test done." severity note;
    WAIT;
  END PROCESS;

	

END TB_ARCH;